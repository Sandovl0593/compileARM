// for Ikarus
// `include "flopenr.v"
// `include "condcheck.v"

module condlogic (
    input wire          clk,
    input wire          reset,
    input wire [3:0]    Cond,
    input wire [3:0]    ALUFlags,
    input wire [1:0]    FlagW,
    input wire          PCS,
    input wire          RegW,
    input wire          MemW,

    output wire         PCSrc,
    output wire         RegWrite,
    output wire         MemWrite
);
    wire [1:0] FlagWrite;
    wire [3:0] Flags;
    wire CondEx;
    flopenr #(2) flagreg1(
        .clk(clk),
        .reset(reset),
        .en(FlagWrite[1]),
        .d(ALUFlags[3:2]),
        .q(Flags[3:2]) // out reg
    );
    flopenr #(2) flagreg0(
        .clk(clk),
        .reset(reset),
        .en(FlagWrite[0]),
        .d(ALUFlags[1:0]),
        .q(Flags[1:0]) // out reg
    );
    condcheck cc(
        .Cond(Cond),
        .Flags(Flags),
        .CondEx(CondEx) // out reg
    );
    assign FlagWrite = FlagW & {2 {CondEx}};
    assign RegWrite = RegW & CondEx;
    assign MemWrite = MemW & CondEx;
    assign PCSrc = PCS & CondEx;
endmodule